------------------------------------------------------------------------------
--  File: alu_tb.vhd
------------------------------------------------------------------------------
--ALU testbench
library IEEE;
use IEEE.std_logic_1164.all;

--Testbench entity is always empty
entity AluTestBench is
end AluTestbench;

architecture Bench of AluTestBench is

 --Component declaration for MUX
component Alu is
	port(
		A_IN, B_IN, C_IN	:	in std_logic_vector(3 downto 0);
		O_OUT				:	out std_logic_vector(3 downto 0));
end component;

--Local signal declarations
--Signal "expected" is not a part of the ALU, it is only used for comparing results.
signal a,b,o,expected	:	std_logic_vector(3 downto 0);
signal c				:	std_logic_vector(1 downto 0);
begin
--Component instantiation of MUX
ALU: Alu port map (a, b, c, o);

--Stimulus process
Stimulus: process
	begin
		--Test F1: Count 1
		c<="00";
		a<="0110";
		b<="0011";
		expected<="0100";
		wait for 3 ns;
		
		a<="1111";
		b<="1111";
		expected<="1000";
		wait for 3 ns;
		
		a<="0000";
		b<="0000";
		expected<="0000";
		wait for 3 ns;

		a<="0110";
		b<="0111";
		expected<="0101";
		wait for 3 ns;
		
		
		
		--Test F2: ROR
		c<="01";
		a<="0110";
		b<="0011";
		expected<="0011";
		wait for 3 ns;
		
		a<="1101";
		b<="1001";
		expected<="1110";
		wait for 3 ns;
		
		a<="0000";
		b<="0110";
		expected<="0000";
		wait for 3 ns;

		a<="1001";
		b<="0111";
		expected<="1100";
		wait for 3 ns;
		
		
		
		--Test F3: set A B 
		c<="10";
		a<="0110";
		b<="0011";
		expected<="1110";
		wait for 3 ns;
		
		a<="1001";
		b<="1010";
		expected<="1101";
		wait for 3 ns;
		
		a<="0000";
		b<="XX10";
		expected<="0100";
		wait for 3 ns;

		a<="1001";
		b<="UU01";
		expected<="1011";
		wait for 3 ns;
		
		
		
		--Test F4: Home TODO
		c<="11";
		a<="0110";
		b<="0011";
		expected<="0000";
		wait for 3 ns;
		
		a<="1111";
		b<="1001";
		expected<="0001";
		wait for 3 ns;
		
		a<="0000";
		b<="0110";
		expected<="0000";
		wait for 3 ns;

		a<="1001";
		b<="0100";
		expected<="0001";
		wait for 3 ns;
		
		wait;  --Suspend
	end process Stimulus;

end Bench;
